# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : sram_1024
#       Words            : 1024
#       Bits             : 32
#       Byte-Write       : 1
#       Aspect Ratio     : 1
#       Output Loading   : 0.5  (pf)
#       Data Slew        : 0.5  (ns)
#       CK Slew          : 0.5  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2022/01/20 01:05:31
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO sram_1024
CLASS BLOCK ;
FOREIGN sram_1024 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 553.040 BY 450.800 ;
SYMMETRY x y r90 ;
SITE core ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 551.920 439.380 553.040 442.620 ;
  LAYER metal3 ;
  RECT 551.920 439.380 553.040 442.620 ;
  LAYER metal2 ;
  RECT 551.920 439.380 553.040 442.620 ;
  LAYER metal1 ;
  RECT 551.920 439.380 553.040 442.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 431.540 553.040 434.780 ;
  LAYER metal3 ;
  RECT 551.920 431.540 553.040 434.780 ;
  LAYER metal2 ;
  RECT 551.920 431.540 553.040 434.780 ;
  LAYER metal1 ;
  RECT 551.920 431.540 553.040 434.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 423.700 553.040 426.940 ;
  LAYER metal3 ;
  RECT 551.920 423.700 553.040 426.940 ;
  LAYER metal2 ;
  RECT 551.920 423.700 553.040 426.940 ;
  LAYER metal1 ;
  RECT 551.920 423.700 553.040 426.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 415.860 553.040 419.100 ;
  LAYER metal3 ;
  RECT 551.920 415.860 553.040 419.100 ;
  LAYER metal2 ;
  RECT 551.920 415.860 553.040 419.100 ;
  LAYER metal1 ;
  RECT 551.920 415.860 553.040 419.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 408.020 553.040 411.260 ;
  LAYER metal3 ;
  RECT 551.920 408.020 553.040 411.260 ;
  LAYER metal2 ;
  RECT 551.920 408.020 553.040 411.260 ;
  LAYER metal1 ;
  RECT 551.920 408.020 553.040 411.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 400.180 553.040 403.420 ;
  LAYER metal3 ;
  RECT 551.920 400.180 553.040 403.420 ;
  LAYER metal2 ;
  RECT 551.920 400.180 553.040 403.420 ;
  LAYER metal1 ;
  RECT 551.920 400.180 553.040 403.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 360.980 553.040 364.220 ;
  LAYER metal3 ;
  RECT 551.920 360.980 553.040 364.220 ;
  LAYER metal2 ;
  RECT 551.920 360.980 553.040 364.220 ;
  LAYER metal1 ;
  RECT 551.920 360.980 553.040 364.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 353.140 553.040 356.380 ;
  LAYER metal3 ;
  RECT 551.920 353.140 553.040 356.380 ;
  LAYER metal2 ;
  RECT 551.920 353.140 553.040 356.380 ;
  LAYER metal1 ;
  RECT 551.920 353.140 553.040 356.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 345.300 553.040 348.540 ;
  LAYER metal3 ;
  RECT 551.920 345.300 553.040 348.540 ;
  LAYER metal2 ;
  RECT 551.920 345.300 553.040 348.540 ;
  LAYER metal1 ;
  RECT 551.920 345.300 553.040 348.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 337.460 553.040 340.700 ;
  LAYER metal3 ;
  RECT 551.920 337.460 553.040 340.700 ;
  LAYER metal2 ;
  RECT 551.920 337.460 553.040 340.700 ;
  LAYER metal1 ;
  RECT 551.920 337.460 553.040 340.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 329.620 553.040 332.860 ;
  LAYER metal3 ;
  RECT 551.920 329.620 553.040 332.860 ;
  LAYER metal2 ;
  RECT 551.920 329.620 553.040 332.860 ;
  LAYER metal1 ;
  RECT 551.920 329.620 553.040 332.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 321.780 553.040 325.020 ;
  LAYER metal3 ;
  RECT 551.920 321.780 553.040 325.020 ;
  LAYER metal2 ;
  RECT 551.920 321.780 553.040 325.020 ;
  LAYER metal1 ;
  RECT 551.920 321.780 553.040 325.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 282.580 553.040 285.820 ;
  LAYER metal3 ;
  RECT 551.920 282.580 553.040 285.820 ;
  LAYER metal2 ;
  RECT 551.920 282.580 553.040 285.820 ;
  LAYER metal1 ;
  RECT 551.920 282.580 553.040 285.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 274.740 553.040 277.980 ;
  LAYER metal3 ;
  RECT 551.920 274.740 553.040 277.980 ;
  LAYER metal2 ;
  RECT 551.920 274.740 553.040 277.980 ;
  LAYER metal1 ;
  RECT 551.920 274.740 553.040 277.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 266.900 553.040 270.140 ;
  LAYER metal3 ;
  RECT 551.920 266.900 553.040 270.140 ;
  LAYER metal2 ;
  RECT 551.920 266.900 553.040 270.140 ;
  LAYER metal1 ;
  RECT 551.920 266.900 553.040 270.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 259.060 553.040 262.300 ;
  LAYER metal3 ;
  RECT 551.920 259.060 553.040 262.300 ;
  LAYER metal2 ;
  RECT 551.920 259.060 553.040 262.300 ;
  LAYER metal1 ;
  RECT 551.920 259.060 553.040 262.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 251.220 553.040 254.460 ;
  LAYER metal3 ;
  RECT 551.920 251.220 553.040 254.460 ;
  LAYER metal2 ;
  RECT 551.920 251.220 553.040 254.460 ;
  LAYER metal1 ;
  RECT 551.920 251.220 553.040 254.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 243.380 553.040 246.620 ;
  LAYER metal3 ;
  RECT 551.920 243.380 553.040 246.620 ;
  LAYER metal2 ;
  RECT 551.920 243.380 553.040 246.620 ;
  LAYER metal1 ;
  RECT 551.920 243.380 553.040 246.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 204.180 553.040 207.420 ;
  LAYER metal3 ;
  RECT 551.920 204.180 553.040 207.420 ;
  LAYER metal2 ;
  RECT 551.920 204.180 553.040 207.420 ;
  LAYER metal1 ;
  RECT 551.920 204.180 553.040 207.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 196.340 553.040 199.580 ;
  LAYER metal3 ;
  RECT 551.920 196.340 553.040 199.580 ;
  LAYER metal2 ;
  RECT 551.920 196.340 553.040 199.580 ;
  LAYER metal1 ;
  RECT 551.920 196.340 553.040 199.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 188.500 553.040 191.740 ;
  LAYER metal3 ;
  RECT 551.920 188.500 553.040 191.740 ;
  LAYER metal2 ;
  RECT 551.920 188.500 553.040 191.740 ;
  LAYER metal1 ;
  RECT 551.920 188.500 553.040 191.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 180.660 553.040 183.900 ;
  LAYER metal3 ;
  RECT 551.920 180.660 553.040 183.900 ;
  LAYER metal2 ;
  RECT 551.920 180.660 553.040 183.900 ;
  LAYER metal1 ;
  RECT 551.920 180.660 553.040 183.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 172.820 553.040 176.060 ;
  LAYER metal3 ;
  RECT 551.920 172.820 553.040 176.060 ;
  LAYER metal2 ;
  RECT 551.920 172.820 553.040 176.060 ;
  LAYER metal1 ;
  RECT 551.920 172.820 553.040 176.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 164.980 553.040 168.220 ;
  LAYER metal3 ;
  RECT 551.920 164.980 553.040 168.220 ;
  LAYER metal2 ;
  RECT 551.920 164.980 553.040 168.220 ;
  LAYER metal1 ;
  RECT 551.920 164.980 553.040 168.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 125.780 553.040 129.020 ;
  LAYER metal3 ;
  RECT 551.920 125.780 553.040 129.020 ;
  LAYER metal2 ;
  RECT 551.920 125.780 553.040 129.020 ;
  LAYER metal1 ;
  RECT 551.920 125.780 553.040 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 117.940 553.040 121.180 ;
  LAYER metal3 ;
  RECT 551.920 117.940 553.040 121.180 ;
  LAYER metal2 ;
  RECT 551.920 117.940 553.040 121.180 ;
  LAYER metal1 ;
  RECT 551.920 117.940 553.040 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 110.100 553.040 113.340 ;
  LAYER metal3 ;
  RECT 551.920 110.100 553.040 113.340 ;
  LAYER metal2 ;
  RECT 551.920 110.100 553.040 113.340 ;
  LAYER metal1 ;
  RECT 551.920 110.100 553.040 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 102.260 553.040 105.500 ;
  LAYER metal3 ;
  RECT 551.920 102.260 553.040 105.500 ;
  LAYER metal2 ;
  RECT 551.920 102.260 553.040 105.500 ;
  LAYER metal1 ;
  RECT 551.920 102.260 553.040 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 94.420 553.040 97.660 ;
  LAYER metal3 ;
  RECT 551.920 94.420 553.040 97.660 ;
  LAYER metal2 ;
  RECT 551.920 94.420 553.040 97.660 ;
  LAYER metal1 ;
  RECT 551.920 94.420 553.040 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 86.580 553.040 89.820 ;
  LAYER metal3 ;
  RECT 551.920 86.580 553.040 89.820 ;
  LAYER metal2 ;
  RECT 551.920 86.580 553.040 89.820 ;
  LAYER metal1 ;
  RECT 551.920 86.580 553.040 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 47.380 553.040 50.620 ;
  LAYER metal3 ;
  RECT 551.920 47.380 553.040 50.620 ;
  LAYER metal2 ;
  RECT 551.920 47.380 553.040 50.620 ;
  LAYER metal1 ;
  RECT 551.920 47.380 553.040 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 39.540 553.040 42.780 ;
  LAYER metal3 ;
  RECT 551.920 39.540 553.040 42.780 ;
  LAYER metal2 ;
  RECT 551.920 39.540 553.040 42.780 ;
  LAYER metal1 ;
  RECT 551.920 39.540 553.040 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 31.700 553.040 34.940 ;
  LAYER metal3 ;
  RECT 551.920 31.700 553.040 34.940 ;
  LAYER metal2 ;
  RECT 551.920 31.700 553.040 34.940 ;
  LAYER metal1 ;
  RECT 551.920 31.700 553.040 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 23.860 553.040 27.100 ;
  LAYER metal3 ;
  RECT 551.920 23.860 553.040 27.100 ;
  LAYER metal2 ;
  RECT 551.920 23.860 553.040 27.100 ;
  LAYER metal1 ;
  RECT 551.920 23.860 553.040 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 16.020 553.040 19.260 ;
  LAYER metal3 ;
  RECT 551.920 16.020 553.040 19.260 ;
  LAYER metal2 ;
  RECT 551.920 16.020 553.040 19.260 ;
  LAYER metal1 ;
  RECT 551.920 16.020 553.040 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 8.180 553.040 11.420 ;
  LAYER metal3 ;
  RECT 551.920 8.180 553.040 11.420 ;
  LAYER metal2 ;
  RECT 551.920 8.180 553.040 11.420 ;
  LAYER metal1 ;
  RECT 551.920 8.180 553.040 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 439.380 1.120 442.620 ;
  LAYER metal3 ;
  RECT 0.000 439.380 1.120 442.620 ;
  LAYER metal2 ;
  RECT 0.000 439.380 1.120 442.620 ;
  LAYER metal1 ;
  RECT 0.000 439.380 1.120 442.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 431.540 1.120 434.780 ;
  LAYER metal3 ;
  RECT 0.000 431.540 1.120 434.780 ;
  LAYER metal2 ;
  RECT 0.000 431.540 1.120 434.780 ;
  LAYER metal1 ;
  RECT 0.000 431.540 1.120 434.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 423.700 1.120 426.940 ;
  LAYER metal3 ;
  RECT 0.000 423.700 1.120 426.940 ;
  LAYER metal2 ;
  RECT 0.000 423.700 1.120 426.940 ;
  LAYER metal1 ;
  RECT 0.000 423.700 1.120 426.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 415.860 1.120 419.100 ;
  LAYER metal3 ;
  RECT 0.000 415.860 1.120 419.100 ;
  LAYER metal2 ;
  RECT 0.000 415.860 1.120 419.100 ;
  LAYER metal1 ;
  RECT 0.000 415.860 1.120 419.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 408.020 1.120 411.260 ;
  LAYER metal3 ;
  RECT 0.000 408.020 1.120 411.260 ;
  LAYER metal2 ;
  RECT 0.000 408.020 1.120 411.260 ;
  LAYER metal1 ;
  RECT 0.000 408.020 1.120 411.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 400.180 1.120 403.420 ;
  LAYER metal3 ;
  RECT 0.000 400.180 1.120 403.420 ;
  LAYER metal2 ;
  RECT 0.000 400.180 1.120 403.420 ;
  LAYER metal1 ;
  RECT 0.000 400.180 1.120 403.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 360.980 1.120 364.220 ;
  LAYER metal3 ;
  RECT 0.000 360.980 1.120 364.220 ;
  LAYER metal2 ;
  RECT 0.000 360.980 1.120 364.220 ;
  LAYER metal1 ;
  RECT 0.000 360.980 1.120 364.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 353.140 1.120 356.380 ;
  LAYER metal3 ;
  RECT 0.000 353.140 1.120 356.380 ;
  LAYER metal2 ;
  RECT 0.000 353.140 1.120 356.380 ;
  LAYER metal1 ;
  RECT 0.000 353.140 1.120 356.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 345.300 1.120 348.540 ;
  LAYER metal3 ;
  RECT 0.000 345.300 1.120 348.540 ;
  LAYER metal2 ;
  RECT 0.000 345.300 1.120 348.540 ;
  LAYER metal1 ;
  RECT 0.000 345.300 1.120 348.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 337.460 1.120 340.700 ;
  LAYER metal3 ;
  RECT 0.000 337.460 1.120 340.700 ;
  LAYER metal2 ;
  RECT 0.000 337.460 1.120 340.700 ;
  LAYER metal1 ;
  RECT 0.000 337.460 1.120 340.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 329.620 1.120 332.860 ;
  LAYER metal3 ;
  RECT 0.000 329.620 1.120 332.860 ;
  LAYER metal2 ;
  RECT 0.000 329.620 1.120 332.860 ;
  LAYER metal1 ;
  RECT 0.000 329.620 1.120 332.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 321.780 1.120 325.020 ;
  LAYER metal3 ;
  RECT 0.000 321.780 1.120 325.020 ;
  LAYER metal2 ;
  RECT 0.000 321.780 1.120 325.020 ;
  LAYER metal1 ;
  RECT 0.000 321.780 1.120 325.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER metal3 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER metal2 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER metal1 ;
  RECT 0.000 282.580 1.120 285.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER metal3 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER metal2 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER metal1 ;
  RECT 0.000 274.740 1.120 277.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER metal3 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER metal2 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER metal1 ;
  RECT 0.000 266.900 1.120 270.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER metal3 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER metal2 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER metal1 ;
  RECT 0.000 259.060 1.120 262.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER metal3 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER metal2 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER metal1 ;
  RECT 0.000 251.220 1.120 254.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER metal3 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER metal2 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER metal1 ;
  RECT 0.000 243.380 1.120 246.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal3 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal2 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal1 ;
  RECT 0.000 204.180 1.120 207.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal3 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal2 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal1 ;
  RECT 0.000 196.340 1.120 199.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal3 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal2 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal1 ;
  RECT 0.000 188.500 1.120 191.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal3 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal2 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal1 ;
  RECT 0.000 180.660 1.120 183.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal3 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal2 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal1 ;
  RECT 0.000 172.820 1.120 176.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal3 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal2 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal1 ;
  RECT 0.000 164.980 1.120 168.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 537.320 449.680 540.860 450.800 ;
  LAYER metal3 ;
  RECT 537.320 449.680 540.860 450.800 ;
  LAYER metal2 ;
  RECT 537.320 449.680 540.860 450.800 ;
  LAYER metal1 ;
  RECT 537.320 449.680 540.860 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 528.640 449.680 532.180 450.800 ;
  LAYER metal3 ;
  RECT 528.640 449.680 532.180 450.800 ;
  LAYER metal2 ;
  RECT 528.640 449.680 532.180 450.800 ;
  LAYER metal1 ;
  RECT 528.640 449.680 532.180 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 485.240 449.680 488.780 450.800 ;
  LAYER metal3 ;
  RECT 485.240 449.680 488.780 450.800 ;
  LAYER metal2 ;
  RECT 485.240 449.680 488.780 450.800 ;
  LAYER metal1 ;
  RECT 485.240 449.680 488.780 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 476.560 449.680 480.100 450.800 ;
  LAYER metal3 ;
  RECT 476.560 449.680 480.100 450.800 ;
  LAYER metal2 ;
  RECT 476.560 449.680 480.100 450.800 ;
  LAYER metal1 ;
  RECT 476.560 449.680 480.100 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 467.880 449.680 471.420 450.800 ;
  LAYER metal3 ;
  RECT 467.880 449.680 471.420 450.800 ;
  LAYER metal2 ;
  RECT 467.880 449.680 471.420 450.800 ;
  LAYER metal1 ;
  RECT 467.880 449.680 471.420 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 459.200 449.680 462.740 450.800 ;
  LAYER metal3 ;
  RECT 459.200 449.680 462.740 450.800 ;
  LAYER metal2 ;
  RECT 459.200 449.680 462.740 450.800 ;
  LAYER metal1 ;
  RECT 459.200 449.680 462.740 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 450.520 449.680 454.060 450.800 ;
  LAYER metal3 ;
  RECT 450.520 449.680 454.060 450.800 ;
  LAYER metal2 ;
  RECT 450.520 449.680 454.060 450.800 ;
  LAYER metal1 ;
  RECT 450.520 449.680 454.060 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 441.840 449.680 445.380 450.800 ;
  LAYER metal3 ;
  RECT 441.840 449.680 445.380 450.800 ;
  LAYER metal2 ;
  RECT 441.840 449.680 445.380 450.800 ;
  LAYER metal1 ;
  RECT 441.840 449.680 445.380 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 398.440 449.680 401.980 450.800 ;
  LAYER metal3 ;
  RECT 398.440 449.680 401.980 450.800 ;
  LAYER metal2 ;
  RECT 398.440 449.680 401.980 450.800 ;
  LAYER metal1 ;
  RECT 398.440 449.680 401.980 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 389.760 449.680 393.300 450.800 ;
  LAYER metal3 ;
  RECT 389.760 449.680 393.300 450.800 ;
  LAYER metal2 ;
  RECT 389.760 449.680 393.300 450.800 ;
  LAYER metal1 ;
  RECT 389.760 449.680 393.300 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 381.080 449.680 384.620 450.800 ;
  LAYER metal3 ;
  RECT 381.080 449.680 384.620 450.800 ;
  LAYER metal2 ;
  RECT 381.080 449.680 384.620 450.800 ;
  LAYER metal1 ;
  RECT 381.080 449.680 384.620 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 372.400 449.680 375.940 450.800 ;
  LAYER metal3 ;
  RECT 372.400 449.680 375.940 450.800 ;
  LAYER metal2 ;
  RECT 372.400 449.680 375.940 450.800 ;
  LAYER metal1 ;
  RECT 372.400 449.680 375.940 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 363.720 449.680 367.260 450.800 ;
  LAYER metal3 ;
  RECT 363.720 449.680 367.260 450.800 ;
  LAYER metal2 ;
  RECT 363.720 449.680 367.260 450.800 ;
  LAYER metal1 ;
  RECT 363.720 449.680 367.260 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 355.040 449.680 358.580 450.800 ;
  LAYER metal3 ;
  RECT 355.040 449.680 358.580 450.800 ;
  LAYER metal2 ;
  RECT 355.040 449.680 358.580 450.800 ;
  LAYER metal1 ;
  RECT 355.040 449.680 358.580 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 311.640 449.680 315.180 450.800 ;
  LAYER metal3 ;
  RECT 311.640 449.680 315.180 450.800 ;
  LAYER metal2 ;
  RECT 311.640 449.680 315.180 450.800 ;
  LAYER metal1 ;
  RECT 311.640 449.680 315.180 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 302.960 449.680 306.500 450.800 ;
  LAYER metal3 ;
  RECT 302.960 449.680 306.500 450.800 ;
  LAYER metal2 ;
  RECT 302.960 449.680 306.500 450.800 ;
  LAYER metal1 ;
  RECT 302.960 449.680 306.500 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 294.280 449.680 297.820 450.800 ;
  LAYER metal3 ;
  RECT 294.280 449.680 297.820 450.800 ;
  LAYER metal2 ;
  RECT 294.280 449.680 297.820 450.800 ;
  LAYER metal1 ;
  RECT 294.280 449.680 297.820 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 285.600 449.680 289.140 450.800 ;
  LAYER metal3 ;
  RECT 285.600 449.680 289.140 450.800 ;
  LAYER metal2 ;
  RECT 285.600 449.680 289.140 450.800 ;
  LAYER metal1 ;
  RECT 285.600 449.680 289.140 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 276.920 449.680 280.460 450.800 ;
  LAYER metal3 ;
  RECT 276.920 449.680 280.460 450.800 ;
  LAYER metal2 ;
  RECT 276.920 449.680 280.460 450.800 ;
  LAYER metal1 ;
  RECT 276.920 449.680 280.460 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 268.240 449.680 271.780 450.800 ;
  LAYER metal3 ;
  RECT 268.240 449.680 271.780 450.800 ;
  LAYER metal2 ;
  RECT 268.240 449.680 271.780 450.800 ;
  LAYER metal1 ;
  RECT 268.240 449.680 271.780 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 224.840 449.680 228.380 450.800 ;
  LAYER metal3 ;
  RECT 224.840 449.680 228.380 450.800 ;
  LAYER metal2 ;
  RECT 224.840 449.680 228.380 450.800 ;
  LAYER metal1 ;
  RECT 224.840 449.680 228.380 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 216.160 449.680 219.700 450.800 ;
  LAYER metal3 ;
  RECT 216.160 449.680 219.700 450.800 ;
  LAYER metal2 ;
  RECT 216.160 449.680 219.700 450.800 ;
  LAYER metal1 ;
  RECT 216.160 449.680 219.700 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 207.480 449.680 211.020 450.800 ;
  LAYER metal3 ;
  RECT 207.480 449.680 211.020 450.800 ;
  LAYER metal2 ;
  RECT 207.480 449.680 211.020 450.800 ;
  LAYER metal1 ;
  RECT 207.480 449.680 211.020 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 198.800 449.680 202.340 450.800 ;
  LAYER metal3 ;
  RECT 198.800 449.680 202.340 450.800 ;
  LAYER metal2 ;
  RECT 198.800 449.680 202.340 450.800 ;
  LAYER metal1 ;
  RECT 198.800 449.680 202.340 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 190.120 449.680 193.660 450.800 ;
  LAYER metal3 ;
  RECT 190.120 449.680 193.660 450.800 ;
  LAYER metal2 ;
  RECT 190.120 449.680 193.660 450.800 ;
  LAYER metal1 ;
  RECT 190.120 449.680 193.660 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 181.440 449.680 184.980 450.800 ;
  LAYER metal3 ;
  RECT 181.440 449.680 184.980 450.800 ;
  LAYER metal2 ;
  RECT 181.440 449.680 184.980 450.800 ;
  LAYER metal1 ;
  RECT 181.440 449.680 184.980 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 138.040 449.680 141.580 450.800 ;
  LAYER metal3 ;
  RECT 138.040 449.680 141.580 450.800 ;
  LAYER metal2 ;
  RECT 138.040 449.680 141.580 450.800 ;
  LAYER metal1 ;
  RECT 138.040 449.680 141.580 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 129.360 449.680 132.900 450.800 ;
  LAYER metal3 ;
  RECT 129.360 449.680 132.900 450.800 ;
  LAYER metal2 ;
  RECT 129.360 449.680 132.900 450.800 ;
  LAYER metal1 ;
  RECT 129.360 449.680 132.900 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 120.680 449.680 124.220 450.800 ;
  LAYER metal3 ;
  RECT 120.680 449.680 124.220 450.800 ;
  LAYER metal2 ;
  RECT 120.680 449.680 124.220 450.800 ;
  LAYER metal1 ;
  RECT 120.680 449.680 124.220 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 112.000 449.680 115.540 450.800 ;
  LAYER metal3 ;
  RECT 112.000 449.680 115.540 450.800 ;
  LAYER metal2 ;
  RECT 112.000 449.680 115.540 450.800 ;
  LAYER metal1 ;
  RECT 112.000 449.680 115.540 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 103.320 449.680 106.860 450.800 ;
  LAYER metal3 ;
  RECT 103.320 449.680 106.860 450.800 ;
  LAYER metal2 ;
  RECT 103.320 449.680 106.860 450.800 ;
  LAYER metal1 ;
  RECT 103.320 449.680 106.860 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 94.640 449.680 98.180 450.800 ;
  LAYER metal3 ;
  RECT 94.640 449.680 98.180 450.800 ;
  LAYER metal2 ;
  RECT 94.640 449.680 98.180 450.800 ;
  LAYER metal1 ;
  RECT 94.640 449.680 98.180 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 51.240 449.680 54.780 450.800 ;
  LAYER metal3 ;
  RECT 51.240 449.680 54.780 450.800 ;
  LAYER metal2 ;
  RECT 51.240 449.680 54.780 450.800 ;
  LAYER metal1 ;
  RECT 51.240 449.680 54.780 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 42.560 449.680 46.100 450.800 ;
  LAYER metal3 ;
  RECT 42.560 449.680 46.100 450.800 ;
  LAYER metal2 ;
  RECT 42.560 449.680 46.100 450.800 ;
  LAYER metal1 ;
  RECT 42.560 449.680 46.100 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 33.880 449.680 37.420 450.800 ;
  LAYER metal3 ;
  RECT 33.880 449.680 37.420 450.800 ;
  LAYER metal2 ;
  RECT 33.880 449.680 37.420 450.800 ;
  LAYER metal1 ;
  RECT 33.880 449.680 37.420 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 25.200 449.680 28.740 450.800 ;
  LAYER metal3 ;
  RECT 25.200 449.680 28.740 450.800 ;
  LAYER metal2 ;
  RECT 25.200 449.680 28.740 450.800 ;
  LAYER metal1 ;
  RECT 25.200 449.680 28.740 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 16.520 449.680 20.060 450.800 ;
  LAYER metal3 ;
  RECT 16.520 449.680 20.060 450.800 ;
  LAYER metal2 ;
  RECT 16.520 449.680 20.060 450.800 ;
  LAYER metal1 ;
  RECT 16.520 449.680 20.060 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 7.840 449.680 11.380 450.800 ;
  LAYER metal3 ;
  RECT 7.840 449.680 11.380 450.800 ;
  LAYER metal2 ;
  RECT 7.840 449.680 11.380 450.800 ;
  LAYER metal1 ;
  RECT 7.840 449.680 11.380 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 541.660 0.000 545.200 1.120 ;
  LAYER metal3 ;
  RECT 541.660 0.000 545.200 1.120 ;
  LAYER metal2 ;
  RECT 541.660 0.000 545.200 1.120 ;
  LAYER metal1 ;
  RECT 541.660 0.000 545.200 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 519.960 0.000 523.500 1.120 ;
  LAYER metal3 ;
  RECT 519.960 0.000 523.500 1.120 ;
  LAYER metal2 ;
  RECT 519.960 0.000 523.500 1.120 ;
  LAYER metal1 ;
  RECT 519.960 0.000 523.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 503.220 0.000 506.760 1.120 ;
  LAYER metal3 ;
  RECT 503.220 0.000 506.760 1.120 ;
  LAYER metal2 ;
  RECT 503.220 0.000 506.760 1.120 ;
  LAYER metal1 ;
  RECT 503.220 0.000 506.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 476.560 0.000 480.100 1.120 ;
  LAYER metal3 ;
  RECT 476.560 0.000 480.100 1.120 ;
  LAYER metal2 ;
  RECT 476.560 0.000 480.100 1.120 ;
  LAYER metal1 ;
  RECT 476.560 0.000 480.100 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 454.860 0.000 458.400 1.120 ;
  LAYER metal3 ;
  RECT 454.860 0.000 458.400 1.120 ;
  LAYER metal2 ;
  RECT 454.860 0.000 458.400 1.120 ;
  LAYER metal1 ;
  RECT 454.860 0.000 458.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER metal3 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER metal2 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER metal1 ;
  RECT 342.020 0.000 345.560 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 320.320 0.000 323.860 1.120 ;
  LAYER metal3 ;
  RECT 320.320 0.000 323.860 1.120 ;
  LAYER metal2 ;
  RECT 320.320 0.000 323.860 1.120 ;
  LAYER metal1 ;
  RECT 320.320 0.000 323.860 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 293.040 0.000 296.580 1.120 ;
  LAYER metal3 ;
  RECT 293.040 0.000 296.580 1.120 ;
  LAYER metal2 ;
  RECT 293.040 0.000 296.580 1.120 ;
  LAYER metal1 ;
  RECT 293.040 0.000 296.580 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 284.360 0.000 287.900 1.120 ;
  LAYER metal3 ;
  RECT 284.360 0.000 287.900 1.120 ;
  LAYER metal2 ;
  RECT 284.360 0.000 287.900 1.120 ;
  LAYER metal1 ;
  RECT 284.360 0.000 287.900 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 257.080 0.000 260.620 1.120 ;
  LAYER metal3 ;
  RECT 257.080 0.000 260.620 1.120 ;
  LAYER metal2 ;
  RECT 257.080 0.000 260.620 1.120 ;
  LAYER metal1 ;
  RECT 257.080 0.000 260.620 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 235.380 0.000 238.920 1.120 ;
  LAYER metal3 ;
  RECT 235.380 0.000 238.920 1.120 ;
  LAYER metal2 ;
  RECT 235.380 0.000 238.920 1.120 ;
  LAYER metal1 ;
  RECT 235.380 0.000 238.920 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal3 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal2 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal1 ;
  RECT 126.880 0.000 130.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER metal3 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER metal2 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER metal1 ;
  RECT 100.220 0.000 103.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER metal3 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER metal2 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER metal1 ;
  RECT 83.480 0.000 87.020 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER metal3 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER metal2 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER metal1 ;
  RECT 56.820 0.000 60.360 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal3 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal2 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal1 ;
  RECT 14.040 0.000 17.580 1.120 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 551.920 435.460 553.040 438.700 ;
  LAYER metal3 ;
  RECT 551.920 435.460 553.040 438.700 ;
  LAYER metal2 ;
  RECT 551.920 435.460 553.040 438.700 ;
  LAYER metal1 ;
  RECT 551.920 435.460 553.040 438.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 427.620 553.040 430.860 ;
  LAYER metal3 ;
  RECT 551.920 427.620 553.040 430.860 ;
  LAYER metal2 ;
  RECT 551.920 427.620 553.040 430.860 ;
  LAYER metal1 ;
  RECT 551.920 427.620 553.040 430.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 419.780 553.040 423.020 ;
  LAYER metal3 ;
  RECT 551.920 419.780 553.040 423.020 ;
  LAYER metal2 ;
  RECT 551.920 419.780 553.040 423.020 ;
  LAYER metal1 ;
  RECT 551.920 419.780 553.040 423.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 411.940 553.040 415.180 ;
  LAYER metal3 ;
  RECT 551.920 411.940 553.040 415.180 ;
  LAYER metal2 ;
  RECT 551.920 411.940 553.040 415.180 ;
  LAYER metal1 ;
  RECT 551.920 411.940 553.040 415.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 404.100 553.040 407.340 ;
  LAYER metal3 ;
  RECT 551.920 404.100 553.040 407.340 ;
  LAYER metal2 ;
  RECT 551.920 404.100 553.040 407.340 ;
  LAYER metal1 ;
  RECT 551.920 404.100 553.040 407.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 364.900 553.040 368.140 ;
  LAYER metal3 ;
  RECT 551.920 364.900 553.040 368.140 ;
  LAYER metal2 ;
  RECT 551.920 364.900 553.040 368.140 ;
  LAYER metal1 ;
  RECT 551.920 364.900 553.040 368.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 357.060 553.040 360.300 ;
  LAYER metal3 ;
  RECT 551.920 357.060 553.040 360.300 ;
  LAYER metal2 ;
  RECT 551.920 357.060 553.040 360.300 ;
  LAYER metal1 ;
  RECT 551.920 357.060 553.040 360.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 349.220 553.040 352.460 ;
  LAYER metal3 ;
  RECT 551.920 349.220 553.040 352.460 ;
  LAYER metal2 ;
  RECT 551.920 349.220 553.040 352.460 ;
  LAYER metal1 ;
  RECT 551.920 349.220 553.040 352.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 341.380 553.040 344.620 ;
  LAYER metal3 ;
  RECT 551.920 341.380 553.040 344.620 ;
  LAYER metal2 ;
  RECT 551.920 341.380 553.040 344.620 ;
  LAYER metal1 ;
  RECT 551.920 341.380 553.040 344.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 333.540 553.040 336.780 ;
  LAYER metal3 ;
  RECT 551.920 333.540 553.040 336.780 ;
  LAYER metal2 ;
  RECT 551.920 333.540 553.040 336.780 ;
  LAYER metal1 ;
  RECT 551.920 333.540 553.040 336.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 325.700 553.040 328.940 ;
  LAYER metal3 ;
  RECT 551.920 325.700 553.040 328.940 ;
  LAYER metal2 ;
  RECT 551.920 325.700 553.040 328.940 ;
  LAYER metal1 ;
  RECT 551.920 325.700 553.040 328.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 286.500 553.040 289.740 ;
  LAYER metal3 ;
  RECT 551.920 286.500 553.040 289.740 ;
  LAYER metal2 ;
  RECT 551.920 286.500 553.040 289.740 ;
  LAYER metal1 ;
  RECT 551.920 286.500 553.040 289.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 278.660 553.040 281.900 ;
  LAYER metal3 ;
  RECT 551.920 278.660 553.040 281.900 ;
  LAYER metal2 ;
  RECT 551.920 278.660 553.040 281.900 ;
  LAYER metal1 ;
  RECT 551.920 278.660 553.040 281.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 270.820 553.040 274.060 ;
  LAYER metal3 ;
  RECT 551.920 270.820 553.040 274.060 ;
  LAYER metal2 ;
  RECT 551.920 270.820 553.040 274.060 ;
  LAYER metal1 ;
  RECT 551.920 270.820 553.040 274.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 262.980 553.040 266.220 ;
  LAYER metal3 ;
  RECT 551.920 262.980 553.040 266.220 ;
  LAYER metal2 ;
  RECT 551.920 262.980 553.040 266.220 ;
  LAYER metal1 ;
  RECT 551.920 262.980 553.040 266.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 255.140 553.040 258.380 ;
  LAYER metal3 ;
  RECT 551.920 255.140 553.040 258.380 ;
  LAYER metal2 ;
  RECT 551.920 255.140 553.040 258.380 ;
  LAYER metal1 ;
  RECT 551.920 255.140 553.040 258.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 247.300 553.040 250.540 ;
  LAYER metal3 ;
  RECT 551.920 247.300 553.040 250.540 ;
  LAYER metal2 ;
  RECT 551.920 247.300 553.040 250.540 ;
  LAYER metal1 ;
  RECT 551.920 247.300 553.040 250.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 208.100 553.040 211.340 ;
  LAYER metal3 ;
  RECT 551.920 208.100 553.040 211.340 ;
  LAYER metal2 ;
  RECT 551.920 208.100 553.040 211.340 ;
  LAYER metal1 ;
  RECT 551.920 208.100 553.040 211.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 200.260 553.040 203.500 ;
  LAYER metal3 ;
  RECT 551.920 200.260 553.040 203.500 ;
  LAYER metal2 ;
  RECT 551.920 200.260 553.040 203.500 ;
  LAYER metal1 ;
  RECT 551.920 200.260 553.040 203.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 192.420 553.040 195.660 ;
  LAYER metal3 ;
  RECT 551.920 192.420 553.040 195.660 ;
  LAYER metal2 ;
  RECT 551.920 192.420 553.040 195.660 ;
  LAYER metal1 ;
  RECT 551.920 192.420 553.040 195.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 184.580 553.040 187.820 ;
  LAYER metal3 ;
  RECT 551.920 184.580 553.040 187.820 ;
  LAYER metal2 ;
  RECT 551.920 184.580 553.040 187.820 ;
  LAYER metal1 ;
  RECT 551.920 184.580 553.040 187.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 176.740 553.040 179.980 ;
  LAYER metal3 ;
  RECT 551.920 176.740 553.040 179.980 ;
  LAYER metal2 ;
  RECT 551.920 176.740 553.040 179.980 ;
  LAYER metal1 ;
  RECT 551.920 176.740 553.040 179.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 168.900 553.040 172.140 ;
  LAYER metal3 ;
  RECT 551.920 168.900 553.040 172.140 ;
  LAYER metal2 ;
  RECT 551.920 168.900 553.040 172.140 ;
  LAYER metal1 ;
  RECT 551.920 168.900 553.040 172.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 129.700 553.040 132.940 ;
  LAYER metal3 ;
  RECT 551.920 129.700 553.040 132.940 ;
  LAYER metal2 ;
  RECT 551.920 129.700 553.040 132.940 ;
  LAYER metal1 ;
  RECT 551.920 129.700 553.040 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 121.860 553.040 125.100 ;
  LAYER metal3 ;
  RECT 551.920 121.860 553.040 125.100 ;
  LAYER metal2 ;
  RECT 551.920 121.860 553.040 125.100 ;
  LAYER metal1 ;
  RECT 551.920 121.860 553.040 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 114.020 553.040 117.260 ;
  LAYER metal3 ;
  RECT 551.920 114.020 553.040 117.260 ;
  LAYER metal2 ;
  RECT 551.920 114.020 553.040 117.260 ;
  LAYER metal1 ;
  RECT 551.920 114.020 553.040 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 106.180 553.040 109.420 ;
  LAYER metal3 ;
  RECT 551.920 106.180 553.040 109.420 ;
  LAYER metal2 ;
  RECT 551.920 106.180 553.040 109.420 ;
  LAYER metal1 ;
  RECT 551.920 106.180 553.040 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 98.340 553.040 101.580 ;
  LAYER metal3 ;
  RECT 551.920 98.340 553.040 101.580 ;
  LAYER metal2 ;
  RECT 551.920 98.340 553.040 101.580 ;
  LAYER metal1 ;
  RECT 551.920 98.340 553.040 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 90.500 553.040 93.740 ;
  LAYER metal3 ;
  RECT 551.920 90.500 553.040 93.740 ;
  LAYER metal2 ;
  RECT 551.920 90.500 553.040 93.740 ;
  LAYER metal1 ;
  RECT 551.920 90.500 553.040 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 51.300 553.040 54.540 ;
  LAYER metal3 ;
  RECT 551.920 51.300 553.040 54.540 ;
  LAYER metal2 ;
  RECT 551.920 51.300 553.040 54.540 ;
  LAYER metal1 ;
  RECT 551.920 51.300 553.040 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 43.460 553.040 46.700 ;
  LAYER metal3 ;
  RECT 551.920 43.460 553.040 46.700 ;
  LAYER metal2 ;
  RECT 551.920 43.460 553.040 46.700 ;
  LAYER metal1 ;
  RECT 551.920 43.460 553.040 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 35.620 553.040 38.860 ;
  LAYER metal3 ;
  RECT 551.920 35.620 553.040 38.860 ;
  LAYER metal2 ;
  RECT 551.920 35.620 553.040 38.860 ;
  LAYER metal1 ;
  RECT 551.920 35.620 553.040 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 27.780 553.040 31.020 ;
  LAYER metal3 ;
  RECT 551.920 27.780 553.040 31.020 ;
  LAYER metal2 ;
  RECT 551.920 27.780 553.040 31.020 ;
  LAYER metal1 ;
  RECT 551.920 27.780 553.040 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 19.940 553.040 23.180 ;
  LAYER metal3 ;
  RECT 551.920 19.940 553.040 23.180 ;
  LAYER metal2 ;
  RECT 551.920 19.940 553.040 23.180 ;
  LAYER metal1 ;
  RECT 551.920 19.940 553.040 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 551.920 12.100 553.040 15.340 ;
  LAYER metal3 ;
  RECT 551.920 12.100 553.040 15.340 ;
  LAYER metal2 ;
  RECT 551.920 12.100 553.040 15.340 ;
  LAYER metal1 ;
  RECT 551.920 12.100 553.040 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 435.460 1.120 438.700 ;
  LAYER metal3 ;
  RECT 0.000 435.460 1.120 438.700 ;
  LAYER metal2 ;
  RECT 0.000 435.460 1.120 438.700 ;
  LAYER metal1 ;
  RECT 0.000 435.460 1.120 438.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 427.620 1.120 430.860 ;
  LAYER metal3 ;
  RECT 0.000 427.620 1.120 430.860 ;
  LAYER metal2 ;
  RECT 0.000 427.620 1.120 430.860 ;
  LAYER metal1 ;
  RECT 0.000 427.620 1.120 430.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 419.780 1.120 423.020 ;
  LAYER metal3 ;
  RECT 0.000 419.780 1.120 423.020 ;
  LAYER metal2 ;
  RECT 0.000 419.780 1.120 423.020 ;
  LAYER metal1 ;
  RECT 0.000 419.780 1.120 423.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 411.940 1.120 415.180 ;
  LAYER metal3 ;
  RECT 0.000 411.940 1.120 415.180 ;
  LAYER metal2 ;
  RECT 0.000 411.940 1.120 415.180 ;
  LAYER metal1 ;
  RECT 0.000 411.940 1.120 415.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 404.100 1.120 407.340 ;
  LAYER metal3 ;
  RECT 0.000 404.100 1.120 407.340 ;
  LAYER metal2 ;
  RECT 0.000 404.100 1.120 407.340 ;
  LAYER metal1 ;
  RECT 0.000 404.100 1.120 407.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 364.900 1.120 368.140 ;
  LAYER metal3 ;
  RECT 0.000 364.900 1.120 368.140 ;
  LAYER metal2 ;
  RECT 0.000 364.900 1.120 368.140 ;
  LAYER metal1 ;
  RECT 0.000 364.900 1.120 368.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 357.060 1.120 360.300 ;
  LAYER metal3 ;
  RECT 0.000 357.060 1.120 360.300 ;
  LAYER metal2 ;
  RECT 0.000 357.060 1.120 360.300 ;
  LAYER metal1 ;
  RECT 0.000 357.060 1.120 360.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 349.220 1.120 352.460 ;
  LAYER metal3 ;
  RECT 0.000 349.220 1.120 352.460 ;
  LAYER metal2 ;
  RECT 0.000 349.220 1.120 352.460 ;
  LAYER metal1 ;
  RECT 0.000 349.220 1.120 352.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 341.380 1.120 344.620 ;
  LAYER metal3 ;
  RECT 0.000 341.380 1.120 344.620 ;
  LAYER metal2 ;
  RECT 0.000 341.380 1.120 344.620 ;
  LAYER metal1 ;
  RECT 0.000 341.380 1.120 344.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 333.540 1.120 336.780 ;
  LAYER metal3 ;
  RECT 0.000 333.540 1.120 336.780 ;
  LAYER metal2 ;
  RECT 0.000 333.540 1.120 336.780 ;
  LAYER metal1 ;
  RECT 0.000 333.540 1.120 336.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 325.700 1.120 328.940 ;
  LAYER metal3 ;
  RECT 0.000 325.700 1.120 328.940 ;
  LAYER metal2 ;
  RECT 0.000 325.700 1.120 328.940 ;
  LAYER metal1 ;
  RECT 0.000 325.700 1.120 328.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 286.500 1.120 289.740 ;
  LAYER metal3 ;
  RECT 0.000 286.500 1.120 289.740 ;
  LAYER metal2 ;
  RECT 0.000 286.500 1.120 289.740 ;
  LAYER metal1 ;
  RECT 0.000 286.500 1.120 289.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER metal3 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER metal2 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER metal1 ;
  RECT 0.000 278.660 1.120 281.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER metal3 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER metal2 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER metal1 ;
  RECT 0.000 270.820 1.120 274.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER metal3 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER metal2 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER metal1 ;
  RECT 0.000 262.980 1.120 266.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER metal3 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER metal2 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER metal1 ;
  RECT 0.000 255.140 1.120 258.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER metal3 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER metal2 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER metal1 ;
  RECT 0.000 247.300 1.120 250.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER metal3 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER metal2 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER metal1 ;
  RECT 0.000 208.100 1.120 211.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal3 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal2 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal1 ;
  RECT 0.000 200.260 1.120 203.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal3 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal2 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal1 ;
  RECT 0.000 192.420 1.120 195.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal3 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal2 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal1 ;
  RECT 0.000 184.580 1.120 187.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal3 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal2 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal1 ;
  RECT 0.000 176.740 1.120 179.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal3 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal2 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal1 ;
  RECT 0.000 168.900 1.120 172.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 541.660 449.680 545.200 450.800 ;
  LAYER metal3 ;
  RECT 541.660 449.680 545.200 450.800 ;
  LAYER metal2 ;
  RECT 541.660 449.680 545.200 450.800 ;
  LAYER metal1 ;
  RECT 541.660 449.680 545.200 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 532.980 449.680 536.520 450.800 ;
  LAYER metal3 ;
  RECT 532.980 449.680 536.520 450.800 ;
  LAYER metal2 ;
  RECT 532.980 449.680 536.520 450.800 ;
  LAYER metal1 ;
  RECT 532.980 449.680 536.520 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 489.580 449.680 493.120 450.800 ;
  LAYER metal3 ;
  RECT 489.580 449.680 493.120 450.800 ;
  LAYER metal2 ;
  RECT 489.580 449.680 493.120 450.800 ;
  LAYER metal1 ;
  RECT 489.580 449.680 493.120 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 480.900 449.680 484.440 450.800 ;
  LAYER metal3 ;
  RECT 480.900 449.680 484.440 450.800 ;
  LAYER metal2 ;
  RECT 480.900 449.680 484.440 450.800 ;
  LAYER metal1 ;
  RECT 480.900 449.680 484.440 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 472.220 449.680 475.760 450.800 ;
  LAYER metal3 ;
  RECT 472.220 449.680 475.760 450.800 ;
  LAYER metal2 ;
  RECT 472.220 449.680 475.760 450.800 ;
  LAYER metal1 ;
  RECT 472.220 449.680 475.760 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 463.540 449.680 467.080 450.800 ;
  LAYER metal3 ;
  RECT 463.540 449.680 467.080 450.800 ;
  LAYER metal2 ;
  RECT 463.540 449.680 467.080 450.800 ;
  LAYER metal1 ;
  RECT 463.540 449.680 467.080 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 454.860 449.680 458.400 450.800 ;
  LAYER metal3 ;
  RECT 454.860 449.680 458.400 450.800 ;
  LAYER metal2 ;
  RECT 454.860 449.680 458.400 450.800 ;
  LAYER metal1 ;
  RECT 454.860 449.680 458.400 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 446.180 449.680 449.720 450.800 ;
  LAYER metal3 ;
  RECT 446.180 449.680 449.720 450.800 ;
  LAYER metal2 ;
  RECT 446.180 449.680 449.720 450.800 ;
  LAYER metal1 ;
  RECT 446.180 449.680 449.720 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 402.780 449.680 406.320 450.800 ;
  LAYER metal3 ;
  RECT 402.780 449.680 406.320 450.800 ;
  LAYER metal2 ;
  RECT 402.780 449.680 406.320 450.800 ;
  LAYER metal1 ;
  RECT 402.780 449.680 406.320 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 394.100 449.680 397.640 450.800 ;
  LAYER metal3 ;
  RECT 394.100 449.680 397.640 450.800 ;
  LAYER metal2 ;
  RECT 394.100 449.680 397.640 450.800 ;
  LAYER metal1 ;
  RECT 394.100 449.680 397.640 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 385.420 449.680 388.960 450.800 ;
  LAYER metal3 ;
  RECT 385.420 449.680 388.960 450.800 ;
  LAYER metal2 ;
  RECT 385.420 449.680 388.960 450.800 ;
  LAYER metal1 ;
  RECT 385.420 449.680 388.960 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 376.740 449.680 380.280 450.800 ;
  LAYER metal3 ;
  RECT 376.740 449.680 380.280 450.800 ;
  LAYER metal2 ;
  RECT 376.740 449.680 380.280 450.800 ;
  LAYER metal1 ;
  RECT 376.740 449.680 380.280 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 368.060 449.680 371.600 450.800 ;
  LAYER metal3 ;
  RECT 368.060 449.680 371.600 450.800 ;
  LAYER metal2 ;
  RECT 368.060 449.680 371.600 450.800 ;
  LAYER metal1 ;
  RECT 368.060 449.680 371.600 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 359.380 449.680 362.920 450.800 ;
  LAYER metal3 ;
  RECT 359.380 449.680 362.920 450.800 ;
  LAYER metal2 ;
  RECT 359.380 449.680 362.920 450.800 ;
  LAYER metal1 ;
  RECT 359.380 449.680 362.920 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.980 449.680 319.520 450.800 ;
  LAYER metal3 ;
  RECT 315.980 449.680 319.520 450.800 ;
  LAYER metal2 ;
  RECT 315.980 449.680 319.520 450.800 ;
  LAYER metal1 ;
  RECT 315.980 449.680 319.520 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 307.300 449.680 310.840 450.800 ;
  LAYER metal3 ;
  RECT 307.300 449.680 310.840 450.800 ;
  LAYER metal2 ;
  RECT 307.300 449.680 310.840 450.800 ;
  LAYER metal1 ;
  RECT 307.300 449.680 310.840 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 298.620 449.680 302.160 450.800 ;
  LAYER metal3 ;
  RECT 298.620 449.680 302.160 450.800 ;
  LAYER metal2 ;
  RECT 298.620 449.680 302.160 450.800 ;
  LAYER metal1 ;
  RECT 298.620 449.680 302.160 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 289.940 449.680 293.480 450.800 ;
  LAYER metal3 ;
  RECT 289.940 449.680 293.480 450.800 ;
  LAYER metal2 ;
  RECT 289.940 449.680 293.480 450.800 ;
  LAYER metal1 ;
  RECT 289.940 449.680 293.480 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 281.260 449.680 284.800 450.800 ;
  LAYER metal3 ;
  RECT 281.260 449.680 284.800 450.800 ;
  LAYER metal2 ;
  RECT 281.260 449.680 284.800 450.800 ;
  LAYER metal1 ;
  RECT 281.260 449.680 284.800 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 272.580 449.680 276.120 450.800 ;
  LAYER metal3 ;
  RECT 272.580 449.680 276.120 450.800 ;
  LAYER metal2 ;
  RECT 272.580 449.680 276.120 450.800 ;
  LAYER metal1 ;
  RECT 272.580 449.680 276.120 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 229.180 449.680 232.720 450.800 ;
  LAYER metal3 ;
  RECT 229.180 449.680 232.720 450.800 ;
  LAYER metal2 ;
  RECT 229.180 449.680 232.720 450.800 ;
  LAYER metal1 ;
  RECT 229.180 449.680 232.720 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 220.500 449.680 224.040 450.800 ;
  LAYER metal3 ;
  RECT 220.500 449.680 224.040 450.800 ;
  LAYER metal2 ;
  RECT 220.500 449.680 224.040 450.800 ;
  LAYER metal1 ;
  RECT 220.500 449.680 224.040 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 211.820 449.680 215.360 450.800 ;
  LAYER metal3 ;
  RECT 211.820 449.680 215.360 450.800 ;
  LAYER metal2 ;
  RECT 211.820 449.680 215.360 450.800 ;
  LAYER metal1 ;
  RECT 211.820 449.680 215.360 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 203.140 449.680 206.680 450.800 ;
  LAYER metal3 ;
  RECT 203.140 449.680 206.680 450.800 ;
  LAYER metal2 ;
  RECT 203.140 449.680 206.680 450.800 ;
  LAYER metal1 ;
  RECT 203.140 449.680 206.680 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 194.460 449.680 198.000 450.800 ;
  LAYER metal3 ;
  RECT 194.460 449.680 198.000 450.800 ;
  LAYER metal2 ;
  RECT 194.460 449.680 198.000 450.800 ;
  LAYER metal1 ;
  RECT 194.460 449.680 198.000 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 185.780 449.680 189.320 450.800 ;
  LAYER metal3 ;
  RECT 185.780 449.680 189.320 450.800 ;
  LAYER metal2 ;
  RECT 185.780 449.680 189.320 450.800 ;
  LAYER metal1 ;
  RECT 185.780 449.680 189.320 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 142.380 449.680 145.920 450.800 ;
  LAYER metal3 ;
  RECT 142.380 449.680 145.920 450.800 ;
  LAYER metal2 ;
  RECT 142.380 449.680 145.920 450.800 ;
  LAYER metal1 ;
  RECT 142.380 449.680 145.920 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 133.700 449.680 137.240 450.800 ;
  LAYER metal3 ;
  RECT 133.700 449.680 137.240 450.800 ;
  LAYER metal2 ;
  RECT 133.700 449.680 137.240 450.800 ;
  LAYER metal1 ;
  RECT 133.700 449.680 137.240 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 125.020 449.680 128.560 450.800 ;
  LAYER metal3 ;
  RECT 125.020 449.680 128.560 450.800 ;
  LAYER metal2 ;
  RECT 125.020 449.680 128.560 450.800 ;
  LAYER metal1 ;
  RECT 125.020 449.680 128.560 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 116.340 449.680 119.880 450.800 ;
  LAYER metal3 ;
  RECT 116.340 449.680 119.880 450.800 ;
  LAYER metal2 ;
  RECT 116.340 449.680 119.880 450.800 ;
  LAYER metal1 ;
  RECT 116.340 449.680 119.880 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 107.660 449.680 111.200 450.800 ;
  LAYER metal3 ;
  RECT 107.660 449.680 111.200 450.800 ;
  LAYER metal2 ;
  RECT 107.660 449.680 111.200 450.800 ;
  LAYER metal1 ;
  RECT 107.660 449.680 111.200 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 98.980 449.680 102.520 450.800 ;
  LAYER metal3 ;
  RECT 98.980 449.680 102.520 450.800 ;
  LAYER metal2 ;
  RECT 98.980 449.680 102.520 450.800 ;
  LAYER metal1 ;
  RECT 98.980 449.680 102.520 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 55.580 449.680 59.120 450.800 ;
  LAYER metal3 ;
  RECT 55.580 449.680 59.120 450.800 ;
  LAYER metal2 ;
  RECT 55.580 449.680 59.120 450.800 ;
  LAYER metal1 ;
  RECT 55.580 449.680 59.120 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 46.900 449.680 50.440 450.800 ;
  LAYER metal3 ;
  RECT 46.900 449.680 50.440 450.800 ;
  LAYER metal2 ;
  RECT 46.900 449.680 50.440 450.800 ;
  LAYER metal1 ;
  RECT 46.900 449.680 50.440 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 38.220 449.680 41.760 450.800 ;
  LAYER metal3 ;
  RECT 38.220 449.680 41.760 450.800 ;
  LAYER metal2 ;
  RECT 38.220 449.680 41.760 450.800 ;
  LAYER metal1 ;
  RECT 38.220 449.680 41.760 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 29.540 449.680 33.080 450.800 ;
  LAYER metal3 ;
  RECT 29.540 449.680 33.080 450.800 ;
  LAYER metal2 ;
  RECT 29.540 449.680 33.080 450.800 ;
  LAYER metal1 ;
  RECT 29.540 449.680 33.080 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 20.860 449.680 24.400 450.800 ;
  LAYER metal3 ;
  RECT 20.860 449.680 24.400 450.800 ;
  LAYER metal2 ;
  RECT 20.860 449.680 24.400 450.800 ;
  LAYER metal1 ;
  RECT 20.860 449.680 24.400 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 12.180 449.680 15.720 450.800 ;
  LAYER metal3 ;
  RECT 12.180 449.680 15.720 450.800 ;
  LAYER metal2 ;
  RECT 12.180 449.680 15.720 450.800 ;
  LAYER metal1 ;
  RECT 12.180 449.680 15.720 450.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 532.980 0.000 536.520 1.120 ;
  LAYER metal3 ;
  RECT 532.980 0.000 536.520 1.120 ;
  LAYER metal2 ;
  RECT 532.980 0.000 536.520 1.120 ;
  LAYER metal1 ;
  RECT 532.980 0.000 536.520 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 511.900 0.000 515.440 1.120 ;
  LAYER metal3 ;
  RECT 511.900 0.000 515.440 1.120 ;
  LAYER metal2 ;
  RECT 511.900 0.000 515.440 1.120 ;
  LAYER metal1 ;
  RECT 511.900 0.000 515.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 490.200 0.000 493.740 1.120 ;
  LAYER metal3 ;
  RECT 490.200 0.000 493.740 1.120 ;
  LAYER metal2 ;
  RECT 490.200 0.000 493.740 1.120 ;
  LAYER metal1 ;
  RECT 490.200 0.000 493.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 463.540 0.000 467.080 1.120 ;
  LAYER metal3 ;
  RECT 463.540 0.000 467.080 1.120 ;
  LAYER metal2 ;
  RECT 463.540 0.000 467.080 1.120 ;
  LAYER metal1 ;
  RECT 463.540 0.000 467.080 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 350.080 0.000 353.620 1.120 ;
  LAYER metal3 ;
  RECT 350.080 0.000 353.620 1.120 ;
  LAYER metal2 ;
  RECT 350.080 0.000 353.620 1.120 ;
  LAYER metal1 ;
  RECT 350.080 0.000 353.620 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 333.960 0.000 337.500 1.120 ;
  LAYER metal3 ;
  RECT 333.960 0.000 337.500 1.120 ;
  LAYER metal2 ;
  RECT 333.960 0.000 337.500 1.120 ;
  LAYER metal1 ;
  RECT 333.960 0.000 337.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER metal3 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER metal2 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER metal1 ;
  RECT 297.380 0.000 300.920 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 288.700 0.000 292.240 1.120 ;
  LAYER metal3 ;
  RECT 288.700 0.000 292.240 1.120 ;
  LAYER metal2 ;
  RECT 288.700 0.000 292.240 1.120 ;
  LAYER metal1 ;
  RECT 288.700 0.000 292.240 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 267.620 0.000 271.160 1.120 ;
  LAYER metal3 ;
  RECT 267.620 0.000 271.160 1.120 ;
  LAYER metal2 ;
  RECT 267.620 0.000 271.160 1.120 ;
  LAYER metal1 ;
  RECT 267.620 0.000 271.160 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 246.540 0.000 250.080 1.120 ;
  LAYER metal3 ;
  RECT 246.540 0.000 250.080 1.120 ;
  LAYER metal2 ;
  RECT 246.540 0.000 250.080 1.120 ;
  LAYER metal1 ;
  RECT 246.540 0.000 250.080 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal3 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal2 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal1 ;
  RECT 139.900 0.000 143.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal3 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal2 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal1 ;
  RECT 113.860 0.000 117.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER metal3 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER metal2 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER metal1 ;
  RECT 92.160 0.000 95.700 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal3 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal2 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal1 ;
  RECT 70.460 0.000 74.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER metal3 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER metal2 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER metal1 ;
  RECT 43.800 0.000 47.340 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END GND
PIN DO31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 539.460 0.000 540.580 1.120 ;
  LAYER metal3 ;
  RECT 539.460 0.000 540.580 1.120 ;
  LAYER metal2 ;
  RECT 539.460 0.000 540.580 1.120 ;
  LAYER metal1 ;
  RECT 539.460 0.000 540.580 1.120 ;
 END
END DO31
PIN DI31
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 530.780 0.000 531.900 1.120 ;
  LAYER metal3 ;
  RECT 530.780 0.000 531.900 1.120 ;
  LAYER metal2 ;
  RECT 530.780 0.000 531.900 1.120 ;
  LAYER metal1 ;
  RECT 530.780 0.000 531.900 1.120 ;
 END
END DI31
PIN DO30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 525.820 0.000 526.940 1.120 ;
  LAYER metal3 ;
  RECT 525.820 0.000 526.940 1.120 ;
  LAYER metal2 ;
  RECT 525.820 0.000 526.940 1.120 ;
  LAYER metal1 ;
  RECT 525.820 0.000 526.940 1.120 ;
 END
END DO30
PIN DI30
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 517.760 0.000 518.880 1.120 ;
  LAYER metal3 ;
  RECT 517.760 0.000 518.880 1.120 ;
  LAYER metal2 ;
  RECT 517.760 0.000 518.880 1.120 ;
  LAYER metal1 ;
  RECT 517.760 0.000 518.880 1.120 ;
 END
END DI30
PIN DO29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 509.700 0.000 510.820 1.120 ;
  LAYER metal3 ;
  RECT 509.700 0.000 510.820 1.120 ;
  LAYER metal2 ;
  RECT 509.700 0.000 510.820 1.120 ;
  LAYER metal1 ;
  RECT 509.700 0.000 510.820 1.120 ;
 END
END DO29
PIN DI29
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 501.020 0.000 502.140 1.120 ;
  LAYER metal3 ;
  RECT 501.020 0.000 502.140 1.120 ;
  LAYER metal2 ;
  RECT 501.020 0.000 502.140 1.120 ;
  LAYER metal1 ;
  RECT 501.020 0.000 502.140 1.120 ;
 END
END DI29
PIN DO28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 496.060 0.000 497.180 1.120 ;
  LAYER metal3 ;
  RECT 496.060 0.000 497.180 1.120 ;
  LAYER metal2 ;
  RECT 496.060 0.000 497.180 1.120 ;
  LAYER metal1 ;
  RECT 496.060 0.000 497.180 1.120 ;
 END
END DO28
PIN DI28
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER metal3 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER metal2 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER metal1 ;
  RECT 488.000 0.000 489.120 1.120 ;
 END
END DI28
PIN DO27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER metal3 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER metal2 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER metal1 ;
  RECT 483.040 0.000 484.160 1.120 ;
 END
END DO27
PIN DI27
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 474.360 0.000 475.480 1.120 ;
  LAYER metal3 ;
  RECT 474.360 0.000 475.480 1.120 ;
  LAYER metal2 ;
  RECT 474.360 0.000 475.480 1.120 ;
  LAYER metal1 ;
  RECT 474.360 0.000 475.480 1.120 ;
 END
END DI27
PIN DO26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER metal3 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER metal2 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER metal1 ;
  RECT 469.400 0.000 470.520 1.120 ;
 END
END DO26
PIN DI26
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 461.340 0.000 462.460 1.120 ;
  LAYER metal3 ;
  RECT 461.340 0.000 462.460 1.120 ;
  LAYER metal2 ;
  RECT 461.340 0.000 462.460 1.120 ;
  LAYER metal1 ;
  RECT 461.340 0.000 462.460 1.120 ;
 END
END DI26
PIN DO25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 452.660 0.000 453.780 1.120 ;
  LAYER metal3 ;
  RECT 452.660 0.000 453.780 1.120 ;
  LAYER metal2 ;
  RECT 452.660 0.000 453.780 1.120 ;
  LAYER metal1 ;
  RECT 452.660 0.000 453.780 1.120 ;
 END
END DO25
PIN DI25
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 444.600 0.000 445.720 1.120 ;
  LAYER metal3 ;
  RECT 444.600 0.000 445.720 1.120 ;
  LAYER metal2 ;
  RECT 444.600 0.000 445.720 1.120 ;
  LAYER metal1 ;
  RECT 444.600 0.000 445.720 1.120 ;
 END
END DI25
PIN DO24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 439.640 0.000 440.760 1.120 ;
  LAYER metal3 ;
  RECT 439.640 0.000 440.760 1.120 ;
  LAYER metal2 ;
  RECT 439.640 0.000 440.760 1.120 ;
  LAYER metal1 ;
  RECT 439.640 0.000 440.760 1.120 ;
 END
END DO24
PIN DI24
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 430.960 0.000 432.080 1.120 ;
  LAYER metal3 ;
  RECT 430.960 0.000 432.080 1.120 ;
  LAYER metal2 ;
  RECT 430.960 0.000 432.080 1.120 ;
  LAYER metal1 ;
  RECT 430.960 0.000 432.080 1.120 ;
 END
END DI24
PIN DO23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 426.620 0.000 427.740 1.120 ;
  LAYER metal3 ;
  RECT 426.620 0.000 427.740 1.120 ;
  LAYER metal2 ;
  RECT 426.620 0.000 427.740 1.120 ;
  LAYER metal1 ;
  RECT 426.620 0.000 427.740 1.120 ;
 END
END DO23
PIN DI23
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 417.940 0.000 419.060 1.120 ;
  LAYER metal3 ;
  RECT 417.940 0.000 419.060 1.120 ;
  LAYER metal2 ;
  RECT 417.940 0.000 419.060 1.120 ;
  LAYER metal1 ;
  RECT 417.940 0.000 419.060 1.120 ;
 END
END DI23
PIN DO22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 412.980 0.000 414.100 1.120 ;
  LAYER metal3 ;
  RECT 412.980 0.000 414.100 1.120 ;
  LAYER metal2 ;
  RECT 412.980 0.000 414.100 1.120 ;
  LAYER metal1 ;
  RECT 412.980 0.000 414.100 1.120 ;
 END
END DO22
PIN DI22
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 404.920 0.000 406.040 1.120 ;
  LAYER metal3 ;
  RECT 404.920 0.000 406.040 1.120 ;
  LAYER metal2 ;
  RECT 404.920 0.000 406.040 1.120 ;
  LAYER metal1 ;
  RECT 404.920 0.000 406.040 1.120 ;
 END
END DI22
PIN DO21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 396.240 0.000 397.360 1.120 ;
  LAYER metal3 ;
  RECT 396.240 0.000 397.360 1.120 ;
  LAYER metal2 ;
  RECT 396.240 0.000 397.360 1.120 ;
  LAYER metal1 ;
  RECT 396.240 0.000 397.360 1.120 ;
 END
END DO21
PIN DI21
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 388.180 0.000 389.300 1.120 ;
  LAYER metal3 ;
  RECT 388.180 0.000 389.300 1.120 ;
  LAYER metal2 ;
  RECT 388.180 0.000 389.300 1.120 ;
  LAYER metal1 ;
  RECT 388.180 0.000 389.300 1.120 ;
 END
END DI21
PIN DO20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 383.220 0.000 384.340 1.120 ;
  LAYER metal3 ;
  RECT 383.220 0.000 384.340 1.120 ;
  LAYER metal2 ;
  RECT 383.220 0.000 384.340 1.120 ;
  LAYER metal1 ;
  RECT 383.220 0.000 384.340 1.120 ;
 END
END DO20
PIN DI20
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 374.540 0.000 375.660 1.120 ;
  LAYER metal3 ;
  RECT 374.540 0.000 375.660 1.120 ;
  LAYER metal2 ;
  RECT 374.540 0.000 375.660 1.120 ;
  LAYER metal1 ;
  RECT 374.540 0.000 375.660 1.120 ;
 END
END DI20
PIN DO19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 369.580 0.000 370.700 1.120 ;
  LAYER metal3 ;
  RECT 369.580 0.000 370.700 1.120 ;
  LAYER metal2 ;
  RECT 369.580 0.000 370.700 1.120 ;
  LAYER metal1 ;
  RECT 369.580 0.000 370.700 1.120 ;
 END
END DO19
PIN DI19
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 361.520 0.000 362.640 1.120 ;
  LAYER metal3 ;
  RECT 361.520 0.000 362.640 1.120 ;
  LAYER metal2 ;
  RECT 361.520 0.000 362.640 1.120 ;
  LAYER metal1 ;
  RECT 361.520 0.000 362.640 1.120 ;
 END
END DI19
PIN DO18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 356.560 0.000 357.680 1.120 ;
  LAYER metal3 ;
  RECT 356.560 0.000 357.680 1.120 ;
  LAYER metal2 ;
  RECT 356.560 0.000 357.680 1.120 ;
  LAYER metal1 ;
  RECT 356.560 0.000 357.680 1.120 ;
 END
END DO18
PIN DI18
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 347.880 0.000 349.000 1.120 ;
  LAYER metal3 ;
  RECT 347.880 0.000 349.000 1.120 ;
  LAYER metal2 ;
  RECT 347.880 0.000 349.000 1.120 ;
  LAYER metal1 ;
  RECT 347.880 0.000 349.000 1.120 ;
 END
END DI18
PIN DO17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 339.820 0.000 340.940 1.120 ;
  LAYER metal3 ;
  RECT 339.820 0.000 340.940 1.120 ;
  LAYER metal2 ;
  RECT 339.820 0.000 340.940 1.120 ;
  LAYER metal1 ;
  RECT 339.820 0.000 340.940 1.120 ;
 END
END DO17
PIN DI17
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 331.760 0.000 332.880 1.120 ;
  LAYER metal3 ;
  RECT 331.760 0.000 332.880 1.120 ;
  LAYER metal2 ;
  RECT 331.760 0.000 332.880 1.120 ;
  LAYER metal1 ;
  RECT 331.760 0.000 332.880 1.120 ;
 END
END DI17
PIN DO16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 326.800 0.000 327.920 1.120 ;
  LAYER metal3 ;
  RECT 326.800 0.000 327.920 1.120 ;
  LAYER metal2 ;
  RECT 326.800 0.000 327.920 1.120 ;
  LAYER metal1 ;
  RECT 326.800 0.000 327.920 1.120 ;
 END
END DO16
PIN DI16
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 318.120 0.000 319.240 1.120 ;
  LAYER metal3 ;
  RECT 318.120 0.000 319.240 1.120 ;
  LAYER metal2 ;
  RECT 318.120 0.000 319.240 1.120 ;
  LAYER metal1 ;
  RECT 318.120 0.000 319.240 1.120 ;
 END
END DI16
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 312.540 0.000 313.660 1.120 ;
  LAYER metal3 ;
  RECT 312.540 0.000 313.660 1.120 ;
  LAYER metal2 ;
  RECT 312.540 0.000 313.660 1.120 ;
  LAYER metal1 ;
  RECT 312.540 0.000 313.660 1.120 ;
 END
END A1
PIN WEB
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 310.680 0.000 311.800 1.120 ;
  LAYER metal3 ;
  RECT 310.680 0.000 311.800 1.120 ;
  LAYER metal2 ;
  RECT 310.680 0.000 311.800 1.120 ;
  LAYER metal1 ;
  RECT 310.680 0.000 311.800 1.120 ;
 END
END WEB
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER metal4 ;
  RECT 305.720 0.000 306.840 1.120 ;
  LAYER metal3 ;
  RECT 305.720 0.000 306.840 1.120 ;
  LAYER metal2 ;
  RECT 305.720 0.000 306.840 1.120 ;
  LAYER metal1 ;
  RECT 305.720 0.000 306.840 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER metal4 ;
  RECT 303.860 0.000 304.980 1.120 ;
  LAYER metal3 ;
  RECT 303.860 0.000 304.980 1.120 ;
  LAYER metal2 ;
  RECT 303.860 0.000 304.980 1.120 ;
  LAYER metal1 ;
  RECT 303.860 0.000 304.980 1.120 ;
 END
END CS
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 282.160 0.000 283.280 1.120 ;
  LAYER metal3 ;
  RECT 282.160 0.000 283.280 1.120 ;
  LAYER metal2 ;
  RECT 282.160 0.000 283.280 1.120 ;
  LAYER metal1 ;
  RECT 282.160 0.000 283.280 1.120 ;
 END
END A2
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER metal4 ;
  RECT 279.060 0.000 280.180 1.120 ;
  LAYER metal3 ;
  RECT 279.060 0.000 280.180 1.120 ;
  LAYER metal2 ;
  RECT 279.060 0.000 280.180 1.120 ;
  LAYER metal1 ;
  RECT 279.060 0.000 280.180 1.120 ;
 END
END CK
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 277.200 0.000 278.320 1.120 ;
  LAYER metal3 ;
  RECT 277.200 0.000 278.320 1.120 ;
  LAYER metal2 ;
  RECT 277.200 0.000 278.320 1.120 ;
  LAYER metal1 ;
  RECT 277.200 0.000 278.320 1.120 ;
 END
END A0
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 272.860 0.000 273.980 1.120 ;
  LAYER metal3 ;
  RECT 272.860 0.000 273.980 1.120 ;
  LAYER metal2 ;
  RECT 272.860 0.000 273.980 1.120 ;
  LAYER metal1 ;
  RECT 272.860 0.000 273.980 1.120 ;
 END
END A3
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 265.420 0.000 266.540 1.120 ;
  LAYER metal3 ;
  RECT 265.420 0.000 266.540 1.120 ;
  LAYER metal2 ;
  RECT 265.420 0.000 266.540 1.120 ;
  LAYER metal1 ;
  RECT 265.420 0.000 266.540 1.120 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 262.320 0.000 263.440 1.120 ;
  LAYER metal3 ;
  RECT 262.320 0.000 263.440 1.120 ;
  LAYER metal2 ;
  RECT 262.320 0.000 263.440 1.120 ;
  LAYER metal1 ;
  RECT 262.320 0.000 263.440 1.120 ;
 END
END A5
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal3 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal2 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal1 ;
  RECT 254.880 0.000 256.000 1.120 ;
 END
END A6
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 251.780 0.000 252.900 1.120 ;
  LAYER metal3 ;
  RECT 251.780 0.000 252.900 1.120 ;
  LAYER metal2 ;
  RECT 251.780 0.000 252.900 1.120 ;
  LAYER metal1 ;
  RECT 251.780 0.000 252.900 1.120 ;
 END
END A7
PIN A8
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 244.340 0.000 245.460 1.120 ;
  LAYER metal3 ;
  RECT 244.340 0.000 245.460 1.120 ;
  LAYER metal2 ;
  RECT 244.340 0.000 245.460 1.120 ;
  LAYER metal1 ;
  RECT 244.340 0.000 245.460 1.120 ;
 END
END A8
PIN A9
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal3 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal2 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal1 ;
  RECT 241.240 0.000 242.360 1.120 ;
 END
END A9
PIN DO15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER metal3 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER metal2 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER metal1 ;
  RECT 233.180 0.000 234.300 1.120 ;
 END
END DO15
PIN DI15
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER metal3 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER metal2 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER metal1 ;
  RECT 224.500 0.000 225.620 1.120 ;
 END
END DI15
PIN DO14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER metal3 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER metal2 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER metal1 ;
  RECT 219.540 0.000 220.660 1.120 ;
 END
END DO14
PIN DI14
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER metal3 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER metal2 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER metal1 ;
  RECT 211.480 0.000 212.600 1.120 ;
 END
END DI14
PIN DO13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER metal3 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER metal2 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER metal1 ;
  RECT 202.800 0.000 203.920 1.120 ;
 END
END DO13
PIN DI13
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER metal3 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER metal2 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER metal1 ;
  RECT 194.740 0.000 195.860 1.120 ;
 END
END DI13
PIN DO12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER metal3 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER metal2 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER metal1 ;
  RECT 189.780 0.000 190.900 1.120 ;
 END
END DO12
PIN DI12
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER metal3 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER metal2 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER metal1 ;
  RECT 181.100 0.000 182.220 1.120 ;
 END
END DI12
PIN DO11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER metal3 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER metal2 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER metal1 ;
  RECT 176.140 0.000 177.260 1.120 ;
 END
END DO11
PIN DI11
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER metal3 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER metal2 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER metal1 ;
  RECT 168.080 0.000 169.200 1.120 ;
 END
END DI11
PIN DO10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER metal3 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER metal2 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER metal1 ;
  RECT 163.120 0.000 164.240 1.120 ;
 END
END DO10
PIN DI10
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER metal3 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER metal2 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER metal1 ;
  RECT 154.440 0.000 155.560 1.120 ;
 END
END DI10
PIN DO9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal3 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal2 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal1 ;
  RECT 146.380 0.000 147.500 1.120 ;
 END
END DO9
PIN DI9
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal3 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal2 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal1 ;
  RECT 137.700 0.000 138.820 1.120 ;
 END
END DI9
PIN DO8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal3 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal2 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal1 ;
  RECT 133.360 0.000 134.480 1.120 ;
 END
END DO8
PIN DI8
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal3 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal2 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal1 ;
  RECT 124.680 0.000 125.800 1.120 ;
 END
END DI8
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER metal3 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER metal2 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER metal1 ;
  RECT 119.720 0.000 120.840 1.120 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER metal3 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER metal2 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER metal1 ;
  RECT 111.660 0.000 112.780 1.120 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER metal3 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER metal2 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER metal1 ;
  RECT 98.020 0.000 99.140 1.120 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER metal3 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER metal2 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER metal1 ;
  RECT 89.960 0.000 91.080 1.120 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER metal3 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER metal2 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER metal1 ;
  RECT 81.280 0.000 82.400 1.120 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER metal3 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER metal2 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER metal1 ;
  RECT 76.320 0.000 77.440 1.120 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER metal3 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER metal2 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER metal1 ;
  RECT 68.260 0.000 69.380 1.120 ;
 END
END DI4
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER metal3 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER metal2 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER metal1 ;
  RECT 63.300 0.000 64.420 1.120 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER metal3 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER metal2 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER metal1 ;
  RECT 54.620 0.000 55.740 1.120 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER metal3 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER metal2 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER metal1 ;
  RECT 50.280 0.000 51.400 1.120 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER metal3 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER metal2 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER metal1 ;
  RECT 41.600 0.000 42.720 1.120 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI0
OBS
  LAYER metal1 SPACING 0.280 ;
  RECT 0.000 0.140 553.040 450.800 ;
  LAYER metal2 SPACING 0.320 ;
  RECT 0.000 0.140 553.040 450.800 ;
  LAYER metal3 SPACING 0.320 ;
  RECT 0.000 0.140 553.040 450.800 ;
  LAYER metal4 SPACING 0.600 ;
  RECT 0.000 0.140 553.040 450.800 ;
  LAYER via ;
  RECT 0.000 0.140 553.040 450.800 ;
  LAYER via2 ;
  RECT 0.000 0.140 553.040 450.800 ;
  LAYER via3 ;
  RECT 0.000 0.140 553.040 450.800 ;
END
END sram_1024
END LIBRARY



